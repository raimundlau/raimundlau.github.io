Common Emitter Amplifier
* A simple common-emitter BJT amplifier circuit
* Input: IN, Output: OUT, Power: VCC, Ground: 0

* Power supply
VCC VCC 0 DC 12V

* Input signal source
VIN IN 0 AC 1V

* Bias resistors
R1 VCC BASE 47k
R2 BASE 0 10k

* Input coupling capacitor
C1 IN BASE 10u

* Transistor
Q1 COLLECTOR BASE EMITTER 2N2222

* Collector resistor
RC VCC COLLECTOR 4.7k

* Emitter resistor
RE EMITTER 0 1k

* Emitter bypass capacitor
CE EMITTER 0 100u

* Output coupling capacitor
C2 COLLECTOR OUT 10u

* Load resistor
RL OUT 0 10k

.END
