RC Low-Pass Filter
* Simple first-order RC low-pass filter

* Input voltage source
V1 INPUT 0 AC 1V

* Filter resistor
R1 INPUT OUTPUT 10k

* Filter capacitor
C1 OUTPUT 0 100n

.END
